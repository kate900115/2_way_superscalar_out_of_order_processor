/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  sys_defs.vh                                         //
//                                                                     //
//  Description :  This file has the macro-defines for macros used in  //
//                 the out of order design.                            //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

`define RS_SIZE 	10
`define PRN_SIZE 	48
`define ROB_SIZE	16
